module Sinv_box_0 (input_data, output_data);
	input [3:0] input_data;
	output reg [3:0] output_data;
	
	always @ (*) begin
		case (input_data)
			4'd0:  output_data = 4'd13;
			4'd1:  output_data = 4'd3;
			4'd2:  output_data = 4'd11;
			4'd3:  output_data = 4'd0;
			4'd4:  output_data = 4'd10;
			4'd5:  output_data = 4'd6;
			4'd6:  output_data = 4'd5;
			4'd7:  output_data = 4'd12;
			4'd8:  output_data = 4'd1;
			4'd9:  output_data = 4'd14;
			4'd10: output_data = 4'd4;
			4'd11: output_data = 4'd7;
			4'd12: output_data = 4'd15;
			4'd13: output_data = 4'd9;
			4'd14: output_data = 4'd8;
			4'd15: output_data = 4'd2;
		endcase
	end
endmodule

module Sinv_box_1 (input_data, output_data);
	input [3:0] input_data;
	output reg [3:0] output_data;
	
	always @ (*) begin
		case (input_data)
			4'd0:  output_data = 4'd5;
			4'd1:  output_data = 4'd8;
			4'd2:  output_data = 4'd2;
			4'd3:  output_data = 4'd14;
			4'd4:  output_data = 4'd15;
			4'd5:  output_data = 4'd6;
			4'd6:  output_data = 4'd12;
			4'd7:  output_data = 4'd3;
			4'd8:  output_data = 4'd11;
			4'd9:  output_data = 4'd4;
			4'd10: output_data = 4'd7;
			4'd11: output_data = 4'd9;
			4'd12: output_data = 4'd1;
			4'd13: output_data = 4'd13;
			4'd14: output_data = 4'd10;
			4'd15: output_data = 4'd0;
		endcase
	end
endmodule

module Sinv_box_2 (input_data, output_data);
	input [3:0] input_data;
	output reg [3:0] output_data;
	
	always @ (*) begin
		case (input_data)
			4'd0:  output_data = 4'd12;
			4'd1:  output_data = 4'd9;
			4'd2:  output_data = 4'd15;
			4'd3:  output_data = 4'd4;
			4'd4:  output_data = 4'd11;
			4'd5:  output_data = 4'd14;
			4'd6:  output_data = 4'd1;
			4'd7:  output_data = 4'd2;
			4'd8:  output_data = 4'd0;
			4'd9:  output_data = 4'd3;
			4'd10: output_data = 4'd6;
			4'd11: output_data = 4'd13;
			4'd12: output_data = 4'd5;
			4'd13: output_data = 4'd8;
			4'd14: output_data = 4'd10;
			4'd15: output_data = 4'd7;
		endcase
	end
endmodule

module Sinv_box_3 (input_data, output_data);
	input [3:0] input_data;
	output reg [3:0] output_data;
	
	always @ (*) begin
		case (input_data)
			4'd0:  output_data = 4'd0;
			4'd1:  output_data = 4'd9;
			4'd2:  output_data = 4'd10;
			4'd3:  output_data = 4'd7;
			4'd4:  output_data = 4'd11;
			4'd5:  output_data = 4'd14;
			4'd6:  output_data = 4'd6;
			4'd7:  output_data = 4'd13;
			4'd8:  output_data = 4'd3;
			4'd9:  output_data = 4'd5;
			4'd10: output_data = 4'd12;
			4'd11: output_data = 4'd2;
			4'd12: output_data = 4'd4;
			4'd13: output_data = 4'd8;
			4'd14: output_data = 4'd15;
			4'd15: output_data = 4'd1;
		endcase
	end
endmodule

module Sinv_box_4 (input_data, output_data);
	input [3:0] input_data;
	output reg [3:0] output_data;
	
	always @ (*) begin
		case (input_data)
			4'd0:  output_data = 4'd5;
			4'd1:  output_data = 4'd0;
			4'd2:  output_data = 4'd8;
			4'd3:  output_data = 4'd3;
			4'd4:  output_data = 4'd10;
			4'd5:  output_data = 4'd9;
			4'd6:  output_data = 4'd7;
			4'd7:  output_data = 4'd14;
			4'd8:  output_data = 4'd2;
			4'd9:  output_data = 4'd12;
			4'd10: output_data = 4'd11;
			4'd11: output_data = 4'd6;
			4'd12: output_data = 4'd4;
			4'd13: output_data = 4'd15;
			4'd14: output_data = 4'd13;
			4'd15: output_data = 4'd1;
		endcase
	end
endmodule

module Sinv_box_5 (input_data, output_data);
	input [3:0] input_data;
	output reg [3:0] output_data;
	
	always @ (*) begin
		case (input_data)
			4'd0:  output_data = 4'd8;
			4'd1:  output_data = 4'd15;
			4'd2:  output_data = 4'd2;
			4'd3:  output_data = 4'd9;
			4'd4:  output_data = 4'd4;
			4'd5:  output_data = 4'd1;
			4'd6:  output_data = 4'd13;
			4'd7:  output_data = 4'd14;
			4'd8:  output_data = 4'd11;
			4'd9:  output_data = 4'd6;
			4'd10: output_data = 4'd5;
			4'd11: output_data = 4'd3;
			4'd12: output_data = 4'd7;
			4'd13: output_data = 4'd12;
			4'd14: output_data = 4'd10;
			4'd15: output_data = 4'd0;
		endcase
	end
endmodule

module Sinv_box_6 (input_data, output_data);
	input [3:0] input_data;
	output reg [3:0] output_data;
	
	always @ (*) begin
		case (input_data)
			4'd0:  output_data = 4'd15;
			4'd1:  output_data = 4'd10;
			4'd2:  output_data = 4'd1;
			4'd3:  output_data = 4'd13;
			4'd4:  output_data = 4'd5;
			4'd5:  output_data = 4'd3;
			4'd6:  output_data = 4'd6;
			4'd7:  output_data = 4'd0;
			4'd8:  output_data = 4'd4;
			4'd9:  output_data = 4'd9;
			4'd10: output_data = 4'd14;
			4'd11: output_data = 4'd7;
			4'd12: output_data = 4'd2;
			4'd13: output_data = 4'd12;
			4'd14: output_data = 4'd8;
			4'd15: output_data = 4'd11;
		endcase
	end
endmodule

module Sinv_box_7 (input_data, output_data);
	input [3:0] input_data;
	output reg [3:0] output_data;
	
	always @ (*) begin
		case (input_data)
			4'd0:  output_data = 4'd3;
			4'd1:  output_data = 4'd0;
			4'd2:  output_data = 4'd6;
			4'd3:  output_data = 4'd13;
			4'd4:  output_data = 4'd9;
			4'd5:  output_data = 4'd14;
			4'd6:  output_data = 4'd15;
			4'd7:  output_data = 4'd8;
			4'd8:  output_data = 4'd5;
			4'd9:  output_data = 4'd12;
			4'd10: output_data = 4'd11;
			4'd11: output_data = 4'd7;
			4'd12: output_data = 4'd10;
			4'd13: output_data = 4'd1;
			4'd14: output_data = 4'd4;
			4'd15: output_data = 4'd2;
		endcase
	end
endmodule